#define
edge , negedge ,posedge edge123
rcmos (rpmos ,rnmos
cmos nmos pmos
supply0 supply1 supply01
tri tri0 tri1 tri01 
triand trior trireg
wand wor wire
scalared vectored scalar vector
inout ,inout (inout
input output
   always@
always 
initial
integer real realtime time reg
highz0 ,highz1 highz01 
(pull0 pull1
strong0 strong1
weak0 weak1 weak
large medium small
parameter
specparam
strong0 strong1
event
parameter
defparam
specparam


#action
assign
deassign
force
release
begin begin :begin )begin
case
casex
casez
function
module
macromodule
primitive
specify
table
task
end
endcase
endfunction
endmodule
endprimitive
endspecify
endtable
endtask
fork
join
default
disable
for
forever
else
ifnone
repeat
wait
while
if if(
and ,and (nand
buf not
bufif0 bufif1 bufif01
notif0 notif1
pulldown pullup
tran tranif0 tranif1
rtran rtranif0 rtranif1
xor nor xnor or