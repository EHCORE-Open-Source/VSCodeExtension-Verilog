#define
always
cmos
defparam
edge
event
highz
highz0
highz1
initial
inout
input
integer
large
medium
negedge
nmos
output
parameter
pmos
posedge
pull0
pull1
rcmos
real
realtime
reg
rnmos
rpmos
scalared
small
specparam
strong
strong0
strong1
supply0
supply1
time
tri
tri0
tri1
triand
trior
trireg
vectored
wand
weak
weak0
weak1
wire
wor

#action
and
assign
begin
buf
bufif0
bufif1
case
casex
casez
deassign
default
disable
else
end
endcase
endfunction
endmodule
endprimitive
endspecify
endtable
endtask
for
force
forever
fork
function
if
ifnone
join
macromodule
module
nand
nor
not
notif0
notif1
or
primitive
pulldown
pullup
release
repeat
rtran
rtranif0
rtranif1
specify
table
task
tran
tranif0
tranif1
wait
while
xnor
xor
